module gcd (clk,
    req_rdy,
    req_val,
    reset,
    resp_rdy,
    resp_val,
    req_msg,
    resp_msg);
 input clk;
 output req_rdy;
 input req_val;
 input reset;
 input resp_rdy;
 output resp_val;
 input [31:0] req_msg;
 output [15:0] resp_msg;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire net17;
 wire net16;
 wire net15;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire net14;
 wire _065_;
 wire _066_;
 wire net13;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire net12;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire net11;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire net10;
 wire _307_;
 wire _308_;
 wire net9;
 wire _310_;
 wire _311_;
 wire net8;
 wire _313_;
 wire _314_;
 wire net7;
 wire _316_;
 wire net6;
 wire net5;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire net4;
 wire _404_;
 wire _405_;
 wire _406_;
 wire net3;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire net2;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire net1;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire _460_;
 wire _461_;
 wire _462_;
 wire _463_;
 wire _464_;
 wire _465_;
 wire _466_;
 wire _467_;
 wire _468_;
 wire _469_;
 wire _470_;
 wire _471_;
 wire _472_;
 wire _473_;
 wire _474_;
 wire _475_;
 wire _476_;
 wire _477_;
 wire _478_;
 wire _479_;
 wire _480_;
 wire _481_;
 wire _482_;
 wire _483_;
 wire _484_;
 wire _485_;
 wire \ctrl.state.out[1] ;
 wire \ctrl.state.out[2] ;
 wire \dpath.a_lt_b$in0[0] ;
 wire \dpath.a_lt_b$in0[10] ;
 wire \dpath.a_lt_b$in0[11] ;
 wire \dpath.a_lt_b$in0[12] ;
 wire \dpath.a_lt_b$in0[13] ;
 wire \dpath.a_lt_b$in0[14] ;
 wire \dpath.a_lt_b$in0[15] ;
 wire \dpath.a_lt_b$in0[1] ;
 wire \dpath.a_lt_b$in0[2] ;
 wire \dpath.a_lt_b$in0[3] ;
 wire \dpath.a_lt_b$in0[4] ;
 wire \dpath.a_lt_b$in0[5] ;
 wire \dpath.a_lt_b$in0[6] ;
 wire \dpath.a_lt_b$in0[7] ;
 wire \dpath.a_lt_b$in0[8] ;
 wire \dpath.a_lt_b$in0[9] ;
 wire \dpath.a_lt_b$in1[0] ;
 wire \dpath.a_lt_b$in1[10] ;
 wire \dpath.a_lt_b$in1[11] ;
 wire \dpath.a_lt_b$in1[12] ;
 wire \dpath.a_lt_b$in1[13] ;
 wire \dpath.a_lt_b$in1[14] ;
 wire \dpath.a_lt_b$in1[15] ;
 wire \dpath.a_lt_b$in1[1] ;
 wire \dpath.a_lt_b$in1[2] ;
 wire \dpath.a_lt_b$in1[3] ;
 wire \dpath.a_lt_b$in1[4] ;
 wire \dpath.a_lt_b$in1[5] ;
 wire \dpath.a_lt_b$in1[6] ;
 wire \dpath.a_lt_b$in1[7] ;
 wire \dpath.a_lt_b$in1[8] ;
 wire \dpath.a_lt_b$in1[9] ;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire clknet_2_0__leaf_clk;
 wire clknet_0_clk;
 wire net56;
 wire net57;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net91;
 wire net110;
 wire net111;
 wire net113;
 wire net114;
 wire net115;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net132;
 wire net133;
 wire net134;
 wire net137;
 wire net138;
 wire net139;
 wire net141;
 wire net143;

 INV_X1 _486_ (.A(net34),
    .ZN(_036_));
 BUF_X1 input17 (.A(req_msg[24]),
    .Z(net17));
 BUF_X1 input16 (.A(req_msg[23]),
    .Z(net16));
 BUF_X1 input15 (.A(req_msg[22]),
    .Z(net15));
 NAND3_X1 _490_ (.A1(_036_),
    .A2(net33),
    .A3(net57),
    .ZN(_040_));
 INV_X2 _491_ (.A(\dpath.a_lt_b$in1[11] ),
    .ZN(_041_));
 INV_X2 _492_ (.A(\dpath.a_lt_b$in1[10] ),
    .ZN(_042_));
 INV_X2 _493_ (.A(\dpath.a_lt_b$in1[9] ),
    .ZN(_043_));
 INV_X2 _494_ (.A(\dpath.a_lt_b$in1[8] ),
    .ZN(_044_));
 NAND4_X1 _495_ (.A1(_041_),
    .A2(_042_),
    .A3(_043_),
    .A4(_044_),
    .ZN(_045_));
 INV_X1 _496_ (.A(\dpath.a_lt_b$in1[15] ),
    .ZN(_046_));
 INV_X2 _497_ (.A(\dpath.a_lt_b$in1[14] ),
    .ZN(_047_));
 INV_X2 _498_ (.A(\dpath.a_lt_b$in1[13] ),
    .ZN(_048_));
 NAND3_X1 _499_ (.A1(_046_),
    .A2(_047_),
    .A3(net59),
    .ZN(_049_));
 NOR3_X1 _500_ (.A1(_045_),
    .A2(net61),
    .A3(_049_),
    .ZN(_050_));
 INV_X2 _501_ (.A(\dpath.a_lt_b$in1[7] ),
    .ZN(_051_));
 INV_X2 _502_ (.A(\dpath.a_lt_b$in1[6] ),
    .ZN(_052_));
 INV_X2 _503_ (.A(\dpath.a_lt_b$in1[5] ),
    .ZN(_053_));
 INV_X2 _504_ (.A(\dpath.a_lt_b$in1[4] ),
    .ZN(_054_));
 NAND4_X1 _505_ (.A1(_051_),
    .A2(_052_),
    .A3(_053_),
    .A4(_054_),
    .ZN(_055_));
 INV_X4 _506_ (.A(\dpath.a_lt_b$in1[3] ),
    .ZN(_056_));
 INV_X2 _507_ (.A(\dpath.a_lt_b$in1[2] ),
    .ZN(_057_));
 INV_X2 _508_ (.A(\dpath.a_lt_b$in1[1] ),
    .ZN(_058_));
 INV_X2 _509_ (.A(\dpath.a_lt_b$in1[0] ),
    .ZN(_059_));
 NAND4_X1 _510_ (.A1(_056_),
    .A2(_057_),
    .A3(_058_),
    .A4(_059_),
    .ZN(_060_));
 NOR2_X1 _511_ (.A1(_055_),
    .A2(_060_),
    .ZN(_061_));
 NAND2_X1 _512_ (.A1(_050_),
    .A2(_061_),
    .ZN(_062_));
 INV_X1 _513_ (.A(_062_),
    .ZN(_063_));
 BUF_X1 input14 (.A(req_msg[21]),
    .Z(net14));
 NAND2_X1 _515_ (.A1(_036_),
    .A2(\ctrl.state.out[2] ),
    .ZN(_065_));
 OAI21_X1 _516_ (.A(_040_),
    .B1(_063_),
    .B2(_065_),
    .ZN(_002_));
 INV_X1 _517_ (.A(\ctrl.state.out[2] ),
    .ZN(_066_));
 BUF_X1 input13 (.A(req_msg[20]),
    .Z(net13));
 AND3_X1 _519_ (.A1(_066_),
    .A2(\ctrl.state.out[1] ),
    .A3(_003_),
    .ZN(net53));
 NAND2_X1 _520_ (.A1(net53),
    .A2(net35),
    .ZN(_068_));
 INV_X1 _521_ (.A(net33),
    .ZN(_069_));
 NAND2_X1 _522_ (.A1(_069_),
    .A2(net57),
    .ZN(_070_));
 NAND3_X1 _523_ (.A1(_068_),
    .A2(_036_),
    .A3(_070_),
    .ZN(_000_));
 NAND3_X1 _524_ (.A1(_068_),
    .A2(_036_),
    .A3(\ctrl.state.out[1] ),
    .ZN(_071_));
 OAI21_X1 _525_ (.A(_071_),
    .B1(_062_),
    .B2(_065_),
    .ZN(_001_));
 INV_X1 _526_ (.A(\dpath.a_lt_b$in0[0] ),
    .ZN(_072_));
 XNOR2_X1 _527_ (.A(_072_),
    .B(\dpath.a_lt_b$in1[0] ),
    .ZN(net37));
 BUF_X1 input12 (.A(req_msg[1]),
    .Z(net12));
 XNOR2_X2 _529_ (.A(\dpath.a_lt_b$in0[1] ),
    .B(\dpath.a_lt_b$in1[1] ),
    .ZN(_074_));
 NOR2_X4 _530_ (.A1(_059_),
    .A2(\dpath.a_lt_b$in0[0] ),
    .ZN(_075_));
 XNOR2_X1 _531_ (.A(net85),
    .B(_075_),
    .ZN(net44));
 NAND2_X2 _532_ (.A1(_058_),
    .A2(\dpath.a_lt_b$in0[1] ),
    .ZN(_076_));
 NOR2_X2 _533_ (.A1(_058_),
    .A2(\dpath.a_lt_b$in0[1] ),
    .ZN(_077_));
 OAI21_X2 _534_ (.A(_076_),
    .B1(_075_),
    .B2(_077_),
    .ZN(_078_));
 NAND2_X2 _535_ (.A1(_057_),
    .A2(\dpath.a_lt_b$in0[2] ),
    .ZN(_079_));
 INV_X1 _536_ (.A(\dpath.a_lt_b$in0[2] ),
    .ZN(_080_));
 NAND2_X4 _537_ (.A1(net65),
    .A2(_080_),
    .ZN(_081_));
 NAND2_X4 _538_ (.A1(_079_),
    .A2(_081_),
    .ZN(_082_));
 XNOR2_X1 _539_ (.A(_078_),
    .B(_082_),
    .ZN(net45));
 INV_X2 _540_ (.A(_075_),
    .ZN(_083_));
 NAND2_X2 _541_ (.A1(_074_),
    .A2(_083_),
    .ZN(_084_));
 NAND2_X1 _542_ (.A1(_076_),
    .A2(_079_),
    .ZN(_085_));
 INV_X1 _543_ (.A(_085_),
    .ZN(_086_));
 NAND2_X4 _544_ (.A1(_084_),
    .A2(_086_),
    .ZN(_087_));
 NAND2_X4 _545_ (.A1(_087_),
    .A2(net139),
    .ZN(_088_));
 XNOR2_X2 _546_ (.A(\dpath.a_lt_b$in1[3] ),
    .B(\dpath.a_lt_b$in0[3] ),
    .ZN(_089_));
 XNOR2_X2 _547_ (.A(_088_),
    .B(net77),
    .ZN(net46));
 NAND2_X4 _548_ (.A1(_056_),
    .A2(\dpath.a_lt_b$in0[3] ),
    .ZN(_090_));
 INV_X2 _549_ (.A(\dpath.a_lt_b$in0[3] ),
    .ZN(_091_));
 NAND2_X4 _550_ (.A1(_091_),
    .A2(net62),
    .ZN(_092_));
 NAND2_X4 _551_ (.A1(_092_),
    .A2(_090_),
    .ZN(_093_));
 NOR2_X4 _552_ (.A1(_093_),
    .A2(_082_),
    .ZN(_094_));
 NAND2_X4 _553_ (.A1(_078_),
    .A2(_094_),
    .ZN(_095_));
 NAND2_X2 _554_ (.A1(_079_),
    .A2(_090_),
    .ZN(_096_));
 NAND2_X4 _555_ (.A1(_092_),
    .A2(_096_),
    .ZN(_097_));
 NAND2_X4 _556_ (.A1(_097_),
    .A2(_095_),
    .ZN(_098_));
 NAND2_X4 _557_ (.A1(_054_),
    .A2(net132),
    .ZN(_099_));
 INV_X1 _558_ (.A(\dpath.a_lt_b$in0[4] ),
    .ZN(_100_));
 NAND2_X2 _559_ (.A1(_100_),
    .A2(\dpath.a_lt_b$in1[4] ),
    .ZN(_101_));
 NAND2_X4 _560_ (.A1(_099_),
    .A2(_101_),
    .ZN(_102_));
 XNOR2_X1 _561_ (.A(net78),
    .B(_102_),
    .ZN(net47));
 INV_X2 _562_ (.A(_090_),
    .ZN(_103_));
 INV_X1 _563_ (.A(_099_),
    .ZN(_104_));
 OAI21_X4 _564_ (.A(net76),
    .B1(_103_),
    .B2(_104_),
    .ZN(_105_));
 INV_X4 _565_ (.A(_102_),
    .ZN(_106_));
 NAND2_X4 _566_ (.A1(_089_),
    .A2(_106_),
    .ZN(_107_));
 OAI21_X4 _567_ (.A(_105_),
    .B1(_088_),
    .B2(net88),
    .ZN(_108_));
 BUF_X1 input11 (.A(req_msg[19]),
    .Z(net11));
 XNOR2_X2 _569_ (.A(\dpath.a_lt_b$in1[5] ),
    .B(\dpath.a_lt_b$in0[5] ),
    .ZN(_110_));
 INV_X1 _570_ (.A(_110_),
    .ZN(_111_));
 XNOR2_X1 _571_ (.A(_108_),
    .B(_111_),
    .ZN(net48));
 NAND2_X1 _572_ (.A1(_053_),
    .A2(\dpath.a_lt_b$in0[5] ),
    .ZN(_112_));
 NAND2_X1 _573_ (.A1(_099_),
    .A2(_112_),
    .ZN(_113_));
 OR2_X2 _574_ (.A1(_053_),
    .A2(\dpath.a_lt_b$in0[5] ),
    .ZN(_114_));
 NAND2_X2 _575_ (.A1(_113_),
    .A2(_114_),
    .ZN(_115_));
 NAND2_X4 _576_ (.A1(_097_),
    .A2(_115_),
    .ZN(_116_));
 INV_X4 _577_ (.A(_116_),
    .ZN(_117_));
 NAND2_X4 _578_ (.A1(_117_),
    .A2(_095_),
    .ZN(_118_));
 NAND2_X1 _579_ (.A1(_106_),
    .A2(_110_),
    .ZN(_119_));
 NAND2_X1 _580_ (.A1(_119_),
    .A2(_115_),
    .ZN(_120_));
 AND2_X4 _581_ (.A1(_118_),
    .A2(_120_),
    .ZN(_121_));
 XNOR2_X2 _582_ (.A(\dpath.a_lt_b$in1[6] ),
    .B(\dpath.a_lt_b$in0[6] ),
    .ZN(_122_));
 INV_X1 _583_ (.A(_122_),
    .ZN(_123_));
 XNOR2_X2 _584_ (.A(net82),
    .B(_123_),
    .ZN(net49));
 NAND2_X4 _585_ (.A1(_110_),
    .A2(_122_),
    .ZN(_124_));
 NOR2_X4 _586_ (.A1(_107_),
    .A2(_124_),
    .ZN(_125_));
 NAND3_X4 _587_ (.A1(_125_),
    .A2(net139),
    .A3(_087_),
    .ZN(_126_));
 NAND2_X1 _588_ (.A1(_052_),
    .A2(net67),
    .ZN(_127_));
 NAND2_X1 _589_ (.A1(_112_),
    .A2(_127_),
    .ZN(_128_));
 INV_X1 _590_ (.A(net67),
    .ZN(_129_));
 NAND2_X1 _591_ (.A1(_129_),
    .A2(net113),
    .ZN(_130_));
 NAND2_X2 _592_ (.A1(_128_),
    .A2(_130_),
    .ZN(_131_));
 OAI21_X2 _593_ (.A(_131_),
    .B1(_105_),
    .B2(_124_),
    .ZN(_132_));
 INV_X2 _594_ (.A(_132_),
    .ZN(_133_));
 NAND2_X4 _595_ (.A1(_126_),
    .A2(_133_),
    .ZN(_134_));
 INV_X1 _596_ (.A(\dpath.a_lt_b$in0[7] ),
    .ZN(_135_));
 NAND2_X1 _597_ (.A1(_051_),
    .A2(_135_),
    .ZN(_136_));
 NAND2_X1 _598_ (.A1(\dpath.a_lt_b$in1[7] ),
    .A2(\dpath.a_lt_b$in0[7] ),
    .ZN(_137_));
 NAND2_X2 _599_ (.A1(_136_),
    .A2(_137_),
    .ZN(_138_));
 INV_X1 _600_ (.A(_138_),
    .ZN(_139_));
 XNOR2_X2 _601_ (.A(_139_),
    .B(net87),
    .ZN(net50));
 NAND2_X2 _602_ (.A1(_122_),
    .A2(_138_),
    .ZN(_140_));
 NOR2_X2 _603_ (.A1(_119_),
    .A2(_140_),
    .ZN(_141_));
 NAND2_X4 _604_ (.A1(_098_),
    .A2(_141_),
    .ZN(_142_));
 NOR2_X2 _605_ (.A1(_140_),
    .A2(_115_),
    .ZN(_143_));
 NAND2_X1 _606_ (.A1(_135_),
    .A2(net115),
    .ZN(_144_));
 INV_X1 _607_ (.A(_127_),
    .ZN(_145_));
 NAND2_X2 _608_ (.A1(_051_),
    .A2(net143),
    .ZN(_146_));
 INV_X2 _609_ (.A(_146_),
    .ZN(_147_));
 OAI21_X4 _610_ (.A(_144_),
    .B1(_145_),
    .B2(_147_),
    .ZN(_148_));
 INV_X2 _611_ (.A(_148_),
    .ZN(_149_));
 NOR2_X4 _612_ (.A1(_143_),
    .A2(_149_),
    .ZN(_150_));
 NAND2_X4 _613_ (.A1(_142_),
    .A2(_150_),
    .ZN(_151_));
 NAND2_X2 _614_ (.A1(_044_),
    .A2(net64),
    .ZN(_152_));
 INV_X1 _615_ (.A(net64),
    .ZN(_153_));
 NAND2_X1 _616_ (.A1(_153_),
    .A2(net72),
    .ZN(_154_));
 NAND2_X1 _617_ (.A1(_152_),
    .A2(_154_),
    .ZN(_155_));
 XNOR2_X2 _618_ (.A(net111),
    .B(_155_),
    .ZN(net51));
 INV_X1 _619_ (.A(_082_),
    .ZN(_156_));
 NAND2_X1 _620_ (.A1(_156_),
    .A2(net85),
    .ZN(_157_));
 NOR2_X2 _621_ (.A1(_157_),
    .A2(net80),
    .ZN(_158_));
 XNOR2_X2 _622_ (.A(\dpath.a_lt_b$in1[8] ),
    .B(\dpath.a_lt_b$in0[8] ),
    .ZN(_159_));
 NAND2_X4 _623_ (.A1(_138_),
    .A2(_159_),
    .ZN(_160_));
 NOR2_X4 _624_ (.A1(_124_),
    .A2(_160_),
    .ZN(_161_));
 NAND3_X2 _625_ (.A1(_158_),
    .A2(_161_),
    .A3(_083_),
    .ZN(_162_));
 NOR2_X1 _626_ (.A1(net81),
    .A2(_102_),
    .ZN(_163_));
 NOR2_X1 _627_ (.A1(_057_),
    .A2(net63),
    .ZN(_164_));
 OAI21_X1 _628_ (.A(_079_),
    .B1(_164_),
    .B2(_076_),
    .ZN(_165_));
 NAND2_X1 _629_ (.A1(_163_),
    .A2(_165_),
    .ZN(_166_));
 NAND2_X1 _630_ (.A1(_166_),
    .A2(_105_),
    .ZN(_167_));
 NAND2_X2 _631_ (.A1(_167_),
    .A2(_161_),
    .ZN(_168_));
 NAND2_X2 _632_ (.A1(_043_),
    .A2(\dpath.a_lt_b$in0[9] ),
    .ZN(_169_));
 INV_X1 _633_ (.A(\dpath.a_lt_b$in0[9] ),
    .ZN(_170_));
 NAND2_X2 _634_ (.A1(_170_),
    .A2(\dpath.a_lt_b$in1[9] ),
    .ZN(_171_));
 NAND2_X4 _635_ (.A1(_169_),
    .A2(_171_),
    .ZN(_172_));
 INV_X4 _636_ (.A(_172_),
    .ZN(_173_));
 NAND2_X1 _637_ (.A1(_146_),
    .A2(_152_),
    .ZN(_174_));
 NAND2_X2 _638_ (.A1(_174_),
    .A2(_154_),
    .ZN(_175_));
 OAI21_X2 _639_ (.A(_175_),
    .B1(_160_),
    .B2(_131_),
    .ZN(_176_));
 INV_X1 _640_ (.A(_176_),
    .ZN(_177_));
 NAND4_X1 _641_ (.A1(_162_),
    .A2(_168_),
    .A3(_173_),
    .A4(_177_),
    .ZN(_178_));
 NAND3_X1 _642_ (.A1(_162_),
    .A2(_168_),
    .A3(_177_),
    .ZN(_179_));
 NAND2_X1 _643_ (.A1(_179_),
    .A2(_172_),
    .ZN(_180_));
 NAND2_X2 _644_ (.A1(_178_),
    .A2(_180_),
    .ZN(net52));
 NAND2_X2 _645_ (.A1(_173_),
    .A2(_159_),
    .ZN(_181_));
 NOR2_X4 _646_ (.A1(_181_),
    .A2(_140_),
    .ZN(_182_));
 NAND3_X2 _647_ (.A1(_118_),
    .A2(_120_),
    .A3(_182_),
    .ZN(_183_));
 NAND2_X1 _648_ (.A1(_152_),
    .A2(_169_),
    .ZN(_184_));
 NAND2_X2 _649_ (.A1(_184_),
    .A2(_171_),
    .ZN(_185_));
 OAI21_X4 _650_ (.A(_185_),
    .B1(_148_),
    .B2(_181_),
    .ZN(_186_));
 INV_X1 _651_ (.A(_186_),
    .ZN(_187_));
 NAND2_X2 _652_ (.A1(_183_),
    .A2(_187_),
    .ZN(_188_));
 NAND2_X4 _653_ (.A1(_042_),
    .A2(net68),
    .ZN(_189_));
 INV_X1 _654_ (.A(\dpath.a_lt_b$in0[10] ),
    .ZN(_190_));
 NAND2_X2 _655_ (.A1(_190_),
    .A2(\dpath.a_lt_b$in1[10] ),
    .ZN(_191_));
 NAND2_X4 _656_ (.A1(_189_),
    .A2(_191_),
    .ZN(_192_));
 NAND2_X2 _657_ (.A1(_188_),
    .A2(_192_),
    .ZN(_193_));
 INV_X1 _658_ (.A(_192_),
    .ZN(_194_));
 NAND3_X1 _659_ (.A1(_183_),
    .A2(_194_),
    .A3(_187_),
    .ZN(_195_));
 NAND2_X2 _660_ (.A1(_193_),
    .A2(_195_),
    .ZN(net38));
 NOR2_X4 _661_ (.A1(_172_),
    .A2(_192_),
    .ZN(_196_));
 INV_X4 _662_ (.A(_196_),
    .ZN(_197_));
 NOR2_X4 _663_ (.A1(_197_),
    .A2(_160_),
    .ZN(_198_));
 NAND2_X1 _664_ (.A1(_132_),
    .A2(_198_),
    .ZN(_199_));
 INV_X1 _665_ (.A(_169_),
    .ZN(_200_));
 INV_X1 _666_ (.A(_189_),
    .ZN(_201_));
 OAI21_X2 _667_ (.A(_191_),
    .B1(_200_),
    .B2(_201_),
    .ZN(_202_));
 OAI21_X4 _668_ (.A(_202_),
    .B1(_197_),
    .B2(_175_),
    .ZN(_203_));
 INV_X1 _669_ (.A(_203_),
    .ZN(_204_));
 NAND2_X1 _670_ (.A1(_199_),
    .A2(_204_),
    .ZN(_205_));
 NAND2_X1 _671_ (.A1(_198_),
    .A2(_125_),
    .ZN(_206_));
 NOR2_X2 _672_ (.A1(_206_),
    .A2(_088_),
    .ZN(_207_));
 NOR2_X1 _673_ (.A1(_205_),
    .A2(_207_),
    .ZN(_208_));
 NAND2_X2 _674_ (.A1(_041_),
    .A2(\dpath.a_lt_b$in0[11] ),
    .ZN(_209_));
 INV_X2 _675_ (.A(\dpath.a_lt_b$in0[11] ),
    .ZN(_210_));
 NAND2_X2 _676_ (.A1(_210_),
    .A2(\dpath.a_lt_b$in1[11] ),
    .ZN(_211_));
 NAND2_X4 _677_ (.A1(_209_),
    .A2(_211_),
    .ZN(_212_));
 NAND2_X1 _678_ (.A1(_208_),
    .A2(_212_),
    .ZN(_213_));
 INV_X4 _679_ (.A(_212_),
    .ZN(_214_));
 OAI21_X1 _680_ (.A(_214_),
    .B1(_205_),
    .B2(_207_),
    .ZN(_215_));
 AND2_X1 _681_ (.A1(_213_),
    .A2(_215_),
    .ZN(net39));
 NOR2_X4 _682_ (.A1(_192_),
    .A2(_212_),
    .ZN(_216_));
 NAND3_X2 _683_ (.A1(_216_),
    .A2(net84),
    .A3(_173_),
    .ZN(_217_));
 INV_X2 _684_ (.A(_217_),
    .ZN(_218_));
 NAND2_X4 _685_ (.A1(_151_),
    .A2(_218_),
    .ZN(_219_));
 INV_X1 _686_ (.A(_185_),
    .ZN(_220_));
 NAND2_X1 _687_ (.A1(_216_),
    .A2(_220_),
    .ZN(_221_));
 INV_X1 _688_ (.A(_209_),
    .ZN(_222_));
 OAI21_X1 _689_ (.A(_211_),
    .B1(_201_),
    .B2(_222_),
    .ZN(_223_));
 NAND2_X1 _690_ (.A1(_221_),
    .A2(_223_),
    .ZN(_224_));
 INV_X1 _691_ (.A(_224_),
    .ZN(_225_));
 NAND2_X4 _692_ (.A1(_219_),
    .A2(_225_),
    .ZN(_226_));
 INV_X2 _693_ (.A(\dpath.a_lt_b$in0[12] ),
    .ZN(_227_));
 NOR2_X4 _694_ (.A1(_227_),
    .A2(\dpath.a_lt_b$in1[12] ),
    .ZN(_228_));
 INV_X2 _695_ (.A(\dpath.a_lt_b$in1[12] ),
    .ZN(_229_));
 NOR2_X4 _696_ (.A1(_229_),
    .A2(\dpath.a_lt_b$in0[12] ),
    .ZN(_230_));
 NOR2_X4 _697_ (.A1(_230_),
    .A2(_228_),
    .ZN(_231_));
 NAND2_X2 _698_ (.A1(_226_),
    .A2(net73),
    .ZN(_232_));
 INV_X1 _699_ (.A(net73),
    .ZN(_233_));
 NAND3_X1 _700_ (.A1(_219_),
    .A2(_233_),
    .A3(_225_),
    .ZN(_234_));
 AND2_X2 _701_ (.A1(_232_),
    .A2(_234_),
    .ZN(net40));
 NAND2_X4 _702_ (.A1(_214_),
    .A2(_231_),
    .ZN(_235_));
 NOR2_X4 _703_ (.A1(_197_),
    .A2(_235_),
    .ZN(_236_));
 AND2_X1 _704_ (.A1(_236_),
    .A2(_161_),
    .ZN(_237_));
 NAND2_X1 _705_ (.A1(_108_),
    .A2(_237_),
    .ZN(_238_));
 NAND2_X1 _706_ (.A1(_176_),
    .A2(_236_),
    .ZN(_239_));
 NOR2_X1 _707_ (.A1(_202_),
    .A2(_235_),
    .ZN(_240_));
 INV_X1 _708_ (.A(_230_),
    .ZN(_241_));
 OAI21_X1 _709_ (.A(_241_),
    .B1(_222_),
    .B2(_228_),
    .ZN(_242_));
 INV_X1 _710_ (.A(_242_),
    .ZN(_243_));
 NOR2_X1 _711_ (.A1(_240_),
    .A2(_243_),
    .ZN(_244_));
 NAND2_X1 _712_ (.A1(_239_),
    .A2(_244_),
    .ZN(_245_));
 INV_X1 _713_ (.A(_245_),
    .ZN(_246_));
 NAND2_X1 _714_ (.A1(_238_),
    .A2(_246_),
    .ZN(_247_));
 INV_X2 _715_ (.A(\dpath.a_lt_b$in0[13] ),
    .ZN(_248_));
 NOR2_X4 _716_ (.A1(_248_),
    .A2(\dpath.a_lt_b$in1[13] ),
    .ZN(_249_));
 NOR2_X4 _717_ (.A1(_048_),
    .A2(\dpath.a_lt_b$in0[13] ),
    .ZN(_250_));
 NOR2_X4 _718_ (.A1(_250_),
    .A2(_249_),
    .ZN(_251_));
 NAND2_X1 _719_ (.A1(_247_),
    .A2(net71),
    .ZN(_252_));
 INV_X1 _720_ (.A(net71),
    .ZN(_253_));
 NAND3_X1 _721_ (.A1(_238_),
    .A2(_253_),
    .A3(_246_),
    .ZN(_254_));
 AND2_X1 _722_ (.A1(_252_),
    .A2(_254_),
    .ZN(net41));
 NAND2_X4 _723_ (.A1(_231_),
    .A2(_251_),
    .ZN(_255_));
 INV_X4 _724_ (.A(_255_),
    .ZN(_256_));
 NAND2_X1 _725_ (.A1(_256_),
    .A2(_216_),
    .ZN(_257_));
 INV_X2 _726_ (.A(_257_),
    .ZN(_258_));
 NAND2_X2 _727_ (.A1(_186_),
    .A2(_258_),
    .ZN(_259_));
 INV_X1 _728_ (.A(_250_),
    .ZN(_260_));
 OAI21_X2 _729_ (.A(_260_),
    .B1(_228_),
    .B2(_249_),
    .ZN(_261_));
 INV_X1 _730_ (.A(_261_),
    .ZN(_262_));
 INV_X1 _731_ (.A(_223_),
    .ZN(_263_));
 AOI21_X2 _732_ (.A(_262_),
    .B1(_263_),
    .B2(_256_),
    .ZN(_264_));
 NAND2_X2 _733_ (.A1(_259_),
    .A2(_264_),
    .ZN(_265_));
 INV_X4 _734_ (.A(_265_),
    .ZN(_266_));
 AND2_X4 _735_ (.A1(_258_),
    .A2(_182_),
    .ZN(_267_));
 NAND2_X4 _736_ (.A1(_121_),
    .A2(_267_),
    .ZN(_268_));
 NAND2_X4 _737_ (.A1(_268_),
    .A2(_266_),
    .ZN(_269_));
 INV_X1 _738_ (.A(\dpath.a_lt_b$in0[14] ),
    .ZN(_270_));
 NOR2_X2 _739_ (.A1(_270_),
    .A2(\dpath.a_lt_b$in1[14] ),
    .ZN(_271_));
 NOR2_X4 _740_ (.A1(_047_),
    .A2(net127),
    .ZN(_272_));
 NOR2_X4 _741_ (.A1(_272_),
    .A2(_271_),
    .ZN(_273_));
 NAND2_X4 _742_ (.A1(_269_),
    .A2(_273_),
    .ZN(_274_));
 INV_X1 _743_ (.A(net128),
    .ZN(_275_));
 NAND3_X2 _744_ (.A1(_266_),
    .A2(_268_),
    .A3(_275_),
    .ZN(_276_));
 AND2_X4 _745_ (.A1(_274_),
    .A2(_276_),
    .ZN(net42));
 NAND2_X2 _746_ (.A1(_251_),
    .A2(_273_),
    .ZN(_277_));
 NOR2_X4 _747_ (.A1(_235_),
    .A2(_277_),
    .ZN(_278_));
 AND2_X2 _748_ (.A1(_198_),
    .A2(_278_),
    .ZN(_279_));
 NAND2_X2 _749_ (.A1(_134_),
    .A2(_279_),
    .ZN(_280_));
 NAND2_X2 _750_ (.A1(_203_),
    .A2(_278_),
    .ZN(_281_));
 INV_X1 _751_ (.A(_271_),
    .ZN(_282_));
 INV_X1 _752_ (.A(net126),
    .ZN(_283_));
 OAI21_X2 _753_ (.A(_282_),
    .B1(_283_),
    .B2(_272_),
    .ZN(_284_));
 INV_X1 _754_ (.A(_277_),
    .ZN(_285_));
 AOI21_X2 _755_ (.A(_284_),
    .B1(_285_),
    .B2(_243_),
    .ZN(_286_));
 NAND2_X2 _756_ (.A1(_281_),
    .A2(_286_),
    .ZN(_287_));
 INV_X2 _757_ (.A(_287_),
    .ZN(_288_));
 NAND2_X2 _758_ (.A1(_280_),
    .A2(_288_),
    .ZN(_289_));
 XNOR2_X1 _759_ (.A(\dpath.a_lt_b$in1[15] ),
    .B(\dpath.a_lt_b$in0[15] ),
    .ZN(_290_));
 NAND2_X2 _760_ (.A1(_289_),
    .A2(_290_),
    .ZN(_291_));
 INV_X1 _761_ (.A(_290_),
    .ZN(_292_));
 NAND3_X1 _762_ (.A1(_280_),
    .A2(_288_),
    .A3(_292_),
    .ZN(_293_));
 AND2_X2 _763_ (.A1(_291_),
    .A2(_293_),
    .ZN(net43));
 NAND2_X1 _764_ (.A1(_273_),
    .A2(_290_),
    .ZN(_294_));
 NOR2_X2 _765_ (.A1(net91),
    .A2(_294_),
    .ZN(_295_));
 AND2_X4 _766_ (.A1(_218_),
    .A2(_295_),
    .ZN(_296_));
 NAND2_X4 _767_ (.A1(net134),
    .A2(_296_),
    .ZN(_297_));
 NAND2_X1 _768_ (.A1(_224_),
    .A2(_295_),
    .ZN(_298_));
 NOR2_X1 _769_ (.A1(_261_),
    .A2(_294_),
    .ZN(_299_));
 NAND2_X1 _770_ (.A1(_046_),
    .A2(\dpath.a_lt_b$in0[15] ),
    .ZN(_300_));
 OAI21_X1 _771_ (.A(_300_),
    .B1(_292_),
    .B2(_282_),
    .ZN(_301_));
 NOR2_X2 _772_ (.A1(_299_),
    .A2(_301_),
    .ZN(_302_));
 NAND2_X2 _773_ (.A1(_298_),
    .A2(_302_),
    .ZN(_303_));
 INV_X4 _774_ (.A(_303_),
    .ZN(_304_));
 NAND2_X4 _775_ (.A1(_304_),
    .A2(_297_),
    .ZN(_305_));
 BUF_X1 input10 (.A(req_msg[18]),
    .Z(net10));
 NAND2_X2 _777_ (.A1(net138),
    .A2(net37),
    .ZN(_307_));
 NAND4_X4 _778_ (.A1(_297_),
    .A2(\ctrl.state.out[2] ),
    .A3(_003_),
    .A4(_304_),
    .ZN(_308_));
 BUF_X1 input9 (.A(req_msg[17]),
    .Z(net9));
 OAI21_X2 _780_ (.A(_307_),
    .B1(net141),
    .B2(_059_),
    .ZN(_310_));
 NOR2_X2 _781_ (.A1(_066_),
    .A2(net57),
    .ZN(_311_));
 BUF_X1 input8 (.A(req_msg[16]),
    .Z(net8));
 NAND2_X1 _783_ (.A1(_310_),
    .A2(_311_),
    .ZN(_313_));
 NOR2_X1 _784_ (.A1(\ctrl.state.out[2] ),
    .A2(net36),
    .ZN(_314_));
 BUF_X1 input7 (.A(req_msg[15]),
    .Z(net7));
 AND2_X1 _786_ (.A1(net56),
    .A2(\dpath.a_lt_b$in0[0] ),
    .ZN(_316_));
 BUF_X1 input6 (.A(req_msg[14]),
    .Z(net6));
 BUF_X1 input5 (.A(req_msg[13]),
    .Z(net5));
 AOI21_X1 _789_ (.A(_316_),
    .B1(net57),
    .B2(net8),
    .ZN(_319_));
 NAND2_X1 _790_ (.A1(_313_),
    .A2(_319_),
    .ZN(_004_));
 NAND2_X2 _791_ (.A1(net137),
    .A2(net138),
    .ZN(_320_));
 OAI21_X2 _792_ (.A(_320_),
    .B1(net141),
    .B2(_042_),
    .ZN(_321_));
 NAND2_X1 _793_ (.A1(_321_),
    .A2(_311_),
    .ZN(_322_));
 AND2_X1 _794_ (.A1(net56),
    .A2(net68),
    .ZN(_323_));
 AOI21_X1 _795_ (.A(_323_),
    .B1(net57),
    .B2(net19),
    .ZN(_324_));
 NAND2_X1 _796_ (.A1(_322_),
    .A2(_324_),
    .ZN(_005_));
 NAND3_X4 _797_ (.A1(_297_),
    .A2(\ctrl.state.out[2] ),
    .A3(_304_),
    .ZN(_325_));
 INV_X4 _798_ (.A(_325_),
    .ZN(_326_));
 NAND3_X1 _799_ (.A1(_326_),
    .A2(net58),
    .A3(_003_),
    .ZN(_327_));
 NAND3_X1 _800_ (.A1(_213_),
    .A2(_215_),
    .A3(net138),
    .ZN(_328_));
 NAND2_X1 _801_ (.A1(_327_),
    .A2(_328_),
    .ZN(_329_));
 NAND2_X1 _802_ (.A1(_329_),
    .A2(_311_),
    .ZN(_330_));
 AND2_X1 _803_ (.A1(_314_),
    .A2(\dpath.a_lt_b$in0[11] ),
    .ZN(_331_));
 AOI21_X1 _804_ (.A(_331_),
    .B1(net36),
    .B2(net20),
    .ZN(_332_));
 NAND2_X1 _805_ (.A1(_330_),
    .A2(_332_),
    .ZN(_006_));
 NAND3_X1 _806_ (.A1(_326_),
    .A2(net60),
    .A3(_003_),
    .ZN(_333_));
 NAND3_X1 _807_ (.A1(net79),
    .A2(_234_),
    .A3(_305_),
    .ZN(_334_));
 NAND2_X1 _808_ (.A1(_333_),
    .A2(_334_),
    .ZN(_335_));
 NAND2_X1 _809_ (.A1(_335_),
    .A2(_311_),
    .ZN(_336_));
 AND2_X1 _810_ (.A1(_314_),
    .A2(\dpath.a_lt_b$in0[12] ),
    .ZN(_337_));
 AOI21_X1 _811_ (.A(_337_),
    .B1(net36),
    .B2(net21),
    .ZN(_338_));
 NAND2_X1 _812_ (.A1(_336_),
    .A2(_338_),
    .ZN(_007_));
 NAND3_X1 _813_ (.A1(_326_),
    .A2(net89),
    .A3(_003_),
    .ZN(_339_));
 NAND3_X1 _814_ (.A1(_252_),
    .A2(_254_),
    .A3(_305_),
    .ZN(_340_));
 NAND2_X1 _815_ (.A1(_339_),
    .A2(_340_),
    .ZN(_341_));
 NAND2_X1 _816_ (.A1(_341_),
    .A2(_311_),
    .ZN(_342_));
 AND2_X1 _817_ (.A1(_314_),
    .A2(\dpath.a_lt_b$in0[13] ),
    .ZN(_343_));
 AOI21_X1 _818_ (.A(_343_),
    .B1(net36),
    .B2(net22),
    .ZN(_344_));
 NAND2_X1 _819_ (.A1(_342_),
    .A2(_344_),
    .ZN(_008_));
 NAND3_X1 _820_ (.A1(_326_),
    .A2(\dpath.a_lt_b$in1[14] ),
    .A3(_003_),
    .ZN(_345_));
 NAND3_X1 _821_ (.A1(net83),
    .A2(_276_),
    .A3(_305_),
    .ZN(_346_));
 NAND2_X1 _822_ (.A1(_345_),
    .A2(_346_),
    .ZN(_347_));
 NAND2_X1 _823_ (.A1(_347_),
    .A2(_311_),
    .ZN(_348_));
 AND2_X1 _824_ (.A1(_314_),
    .A2(\dpath.a_lt_b$in0[14] ),
    .ZN(_349_));
 AOI21_X1 _825_ (.A(_349_),
    .B1(net36),
    .B2(net24),
    .ZN(_350_));
 NAND2_X1 _826_ (.A1(_348_),
    .A2(_350_),
    .ZN(_009_));
 NAND3_X1 _827_ (.A1(_326_),
    .A2(\dpath.a_lt_b$in1[15] ),
    .A3(_003_),
    .ZN(_351_));
 NAND3_X1 _828_ (.A1(_291_),
    .A2(_293_),
    .A3(_305_),
    .ZN(_352_));
 NAND2_X1 _829_ (.A1(_351_),
    .A2(_352_),
    .ZN(_353_));
 NAND2_X1 _830_ (.A1(_353_),
    .A2(_311_),
    .ZN(_354_));
 AND2_X1 _831_ (.A1(_314_),
    .A2(\dpath.a_lt_b$in0[15] ),
    .ZN(_355_));
 AOI21_X1 _832_ (.A(_355_),
    .B1(net36),
    .B2(net25),
    .ZN(_356_));
 NAND2_X1 _833_ (.A1(_354_),
    .A2(_356_),
    .ZN(_010_));
 NAND2_X2 _834_ (.A1(net138),
    .A2(net44),
    .ZN(_357_));
 OAI21_X2 _835_ (.A(_357_),
    .B1(_308_),
    .B2(_058_),
    .ZN(_358_));
 NAND2_X1 _836_ (.A1(_358_),
    .A2(_311_),
    .ZN(_359_));
 AND2_X1 _837_ (.A1(net56),
    .A2(\dpath.a_lt_b$in0[1] ),
    .ZN(_360_));
 AOI21_X1 _838_ (.A(_360_),
    .B1(net57),
    .B2(net9),
    .ZN(_361_));
 NAND2_X1 _839_ (.A1(_359_),
    .A2(_361_),
    .ZN(_011_));
 NAND2_X2 _840_ (.A1(net138),
    .A2(net45),
    .ZN(_362_));
 OAI21_X2 _841_ (.A(_362_),
    .B1(_308_),
    .B2(_057_),
    .ZN(_363_));
 NAND2_X1 _842_ (.A1(_363_),
    .A2(_311_),
    .ZN(_364_));
 AND2_X1 _843_ (.A1(net56),
    .A2(\dpath.a_lt_b$in0[2] ),
    .ZN(_365_));
 AOI21_X1 _844_ (.A(_365_),
    .B1(net57),
    .B2(net10),
    .ZN(_366_));
 NAND2_X1 _845_ (.A1(_364_),
    .A2(_366_),
    .ZN(_012_));
 NAND2_X2 _846_ (.A1(_305_),
    .A2(net46),
    .ZN(_367_));
 OAI21_X2 _847_ (.A(_367_),
    .B1(_056_),
    .B2(_308_),
    .ZN(_368_));
 NAND2_X1 _848_ (.A1(_368_),
    .A2(_311_),
    .ZN(_369_));
 AND2_X1 _849_ (.A1(net56),
    .A2(\dpath.a_lt_b$in0[3] ),
    .ZN(_370_));
 AOI21_X1 _850_ (.A(_370_),
    .B1(net57),
    .B2(net11),
    .ZN(_371_));
 NAND2_X1 _851_ (.A1(_371_),
    .A2(_369_),
    .ZN(_013_));
 NAND2_X2 _852_ (.A1(net138),
    .A2(net47),
    .ZN(_372_));
 OAI21_X2 _853_ (.A(_372_),
    .B1(net141),
    .B2(_054_),
    .ZN(_373_));
 NAND2_X1 _854_ (.A1(_373_),
    .A2(_311_),
    .ZN(_374_));
 AND2_X1 _855_ (.A1(net56),
    .A2(net75),
    .ZN(_375_));
 AOI21_X1 _856_ (.A(_375_),
    .B1(net57),
    .B2(net13),
    .ZN(_376_));
 NAND2_X1 _857_ (.A1(_374_),
    .A2(_376_),
    .ZN(_014_));
 NAND2_X2 _858_ (.A1(net48),
    .A2(_305_),
    .ZN(_377_));
 OAI21_X2 _859_ (.A(_377_),
    .B1(net141),
    .B2(_053_),
    .ZN(_378_));
 NAND2_X1 _860_ (.A1(_378_),
    .A2(_311_),
    .ZN(_379_));
 AND2_X1 _861_ (.A1(net56),
    .A2(net66),
    .ZN(_380_));
 AOI21_X1 _862_ (.A(_380_),
    .B1(net57),
    .B2(net14),
    .ZN(_381_));
 NAND2_X1 _863_ (.A1(_379_),
    .A2(_381_),
    .ZN(_015_));
 NAND2_X2 _864_ (.A1(net49),
    .A2(net138),
    .ZN(_382_));
 OAI21_X2 _865_ (.A(_382_),
    .B1(net141),
    .B2(_052_),
    .ZN(_383_));
 NAND2_X1 _866_ (.A1(_383_),
    .A2(_311_),
    .ZN(_384_));
 AND2_X1 _867_ (.A1(net56),
    .A2(net67),
    .ZN(_385_));
 AOI21_X1 _868_ (.A(_385_),
    .B1(net57),
    .B2(net15),
    .ZN(_386_));
 NAND2_X1 _869_ (.A1(_384_),
    .A2(_386_),
    .ZN(_016_));
 NAND2_X2 _870_ (.A1(net133),
    .A2(_305_),
    .ZN(_387_));
 OAI21_X2 _871_ (.A(_387_),
    .B1(_308_),
    .B2(_051_),
    .ZN(_388_));
 NAND2_X1 _872_ (.A1(_388_),
    .A2(_311_),
    .ZN(_389_));
 AND2_X1 _873_ (.A1(net56),
    .A2(net143),
    .ZN(_390_));
 AOI21_X1 _874_ (.A(_390_),
    .B1(net57),
    .B2(net16),
    .ZN(_391_));
 NAND2_X1 _875_ (.A1(_389_),
    .A2(_391_),
    .ZN(_017_));
 NAND2_X2 _876_ (.A1(net110),
    .A2(net138),
    .ZN(_392_));
 OAI21_X2 _877_ (.A(_392_),
    .B1(_308_),
    .B2(_044_),
    .ZN(_393_));
 NAND2_X1 _878_ (.A1(_393_),
    .A2(_311_),
    .ZN(_394_));
 AND2_X1 _879_ (.A1(net56),
    .A2(\dpath.a_lt_b$in0[8] ),
    .ZN(_395_));
 AOI21_X1 _880_ (.A(_395_),
    .B1(net36),
    .B2(net17),
    .ZN(_396_));
 NAND2_X1 _881_ (.A1(_394_),
    .A2(_396_),
    .ZN(_018_));
 NAND2_X1 _882_ (.A1(net52),
    .A2(_305_),
    .ZN(_397_));
 OAI21_X2 _883_ (.A(_397_),
    .B1(_308_),
    .B2(_043_),
    .ZN(_398_));
 NAND2_X1 _884_ (.A1(_398_),
    .A2(_311_),
    .ZN(_399_));
 AND2_X1 _885_ (.A1(net56),
    .A2(\dpath.a_lt_b$in0[9] ),
    .ZN(_400_));
 AOI21_X1 _886_ (.A(_400_),
    .B1(net36),
    .B2(net18),
    .ZN(_401_));
 NAND2_X1 _887_ (.A1(_399_),
    .A2(_401_),
    .ZN(_019_));
 NAND2_X4 _888_ (.A1(_325_),
    .A2(_003_),
    .ZN(_402_));
 BUF_X1 input4 (.A(req_msg[12]),
    .Z(net4));
 NAND2_X1 _890_ (.A1(net57),
    .A2(net1),
    .ZN(_404_));
 OAI21_X1 _891_ (.A(_404_),
    .B1(_072_),
    .B2(net57),
    .ZN(_405_));
 NAND2_X1 _892_ (.A1(_402_),
    .A2(_405_),
    .ZN(_406_));
 BUF_X1 input3 (.A(req_msg[11]),
    .Z(net3));
 OAI21_X1 _894_ (.A(_406_),
    .B1(_059_),
    .B2(_402_),
    .ZN(_020_));
 NAND2_X1 _895_ (.A1(net57),
    .A2(net2),
    .ZN(_408_));
 OAI21_X1 _896_ (.A(_408_),
    .B1(_190_),
    .B2(net57),
    .ZN(_409_));
 NAND2_X1 _897_ (.A1(_402_),
    .A2(_409_),
    .ZN(_410_));
 OAI21_X1 _898_ (.A(_410_),
    .B1(_042_),
    .B2(_402_),
    .ZN(_021_));
 NAND2_X1 _899_ (.A1(net36),
    .A2(net3),
    .ZN(_411_));
 BUF_X1 input2 (.A(req_msg[10]),
    .Z(net2));
 OAI21_X1 _901_ (.A(_411_),
    .B1(_210_),
    .B2(net36),
    .ZN(_413_));
 NAND2_X1 _902_ (.A1(_402_),
    .A2(_413_),
    .ZN(_414_));
 OAI21_X1 _903_ (.A(_414_),
    .B1(_041_),
    .B2(_402_),
    .ZN(_022_));
 NAND2_X1 _904_ (.A1(net36),
    .A2(net4),
    .ZN(_415_));
 OAI21_X1 _905_ (.A(_415_),
    .B1(net86),
    .B2(net36),
    .ZN(_416_));
 NAND2_X1 _906_ (.A1(_402_),
    .A2(_416_),
    .ZN(_417_));
 OAI21_X1 _907_ (.A(_417_),
    .B1(_229_),
    .B2(_402_),
    .ZN(_023_));
 BUF_X1 input1 (.A(req_msg[0]),
    .Z(net1));
 NAND2_X1 _909_ (.A1(net36),
    .A2(net5),
    .ZN(_419_));
 OAI21_X1 _910_ (.A(_419_),
    .B1(net70),
    .B2(net36),
    .ZN(_420_));
 NAND2_X1 _911_ (.A1(_402_),
    .A2(_420_),
    .ZN(_421_));
 OAI21_X1 _912_ (.A(_421_),
    .B1(net59),
    .B2(_402_),
    .ZN(_024_));
 NAND2_X1 _913_ (.A1(net36),
    .A2(net6),
    .ZN(_422_));
 OAI21_X1 _914_ (.A(_422_),
    .B1(_270_),
    .B2(net36),
    .ZN(_423_));
 NAND2_X1 _915_ (.A1(_402_),
    .A2(_423_),
    .ZN(_424_));
 OAI21_X1 _916_ (.A(_424_),
    .B1(_047_),
    .B2(_402_),
    .ZN(_025_));
 MUX2_X1 _917_ (.A(\dpath.a_lt_b$in0[15] ),
    .B(net7),
    .S(net36),
    .Z(_425_));
 NAND2_X1 _918_ (.A1(_402_),
    .A2(_425_),
    .ZN(_426_));
 OAI21_X1 _919_ (.A(_426_),
    .B1(_046_),
    .B2(_402_),
    .ZN(_026_));
 MUX2_X1 _920_ (.A(\dpath.a_lt_b$in0[1] ),
    .B(net12),
    .S(net57),
    .Z(_427_));
 NAND2_X1 _921_ (.A1(_402_),
    .A2(_427_),
    .ZN(_428_));
 OAI21_X1 _922_ (.A(_428_),
    .B1(_058_),
    .B2(_402_),
    .ZN(_027_));
 NAND2_X1 _923_ (.A1(net57),
    .A2(net23),
    .ZN(_429_));
 OAI21_X1 _924_ (.A(_429_),
    .B1(_080_),
    .B2(net57),
    .ZN(_430_));
 NAND2_X1 _925_ (.A1(_402_),
    .A2(_430_),
    .ZN(_431_));
 OAI21_X1 _926_ (.A(_431_),
    .B1(_057_),
    .B2(_402_),
    .ZN(_028_));
 NAND2_X1 _927_ (.A1(net57),
    .A2(net26),
    .ZN(_432_));
 OAI21_X1 _928_ (.A(_432_),
    .B1(net69),
    .B2(net57),
    .ZN(_433_));
 NAND2_X1 _929_ (.A1(_402_),
    .A2(_433_),
    .ZN(_434_));
 OAI21_X1 _930_ (.A(_434_),
    .B1(_056_),
    .B2(_402_),
    .ZN(_029_));
 NAND2_X1 _931_ (.A1(net57),
    .A2(net27),
    .ZN(_435_));
 OAI21_X1 _932_ (.A(_435_),
    .B1(_100_),
    .B2(net57),
    .ZN(_436_));
 NAND2_X1 _933_ (.A1(_402_),
    .A2(_436_),
    .ZN(_437_));
 OAI21_X1 _934_ (.A(_437_),
    .B1(_054_),
    .B2(_402_),
    .ZN(_030_));
 MUX2_X1 _935_ (.A(net66),
    .B(net28),
    .S(net57),
    .Z(_438_));
 NAND2_X1 _936_ (.A1(_402_),
    .A2(_438_),
    .ZN(_439_));
 OAI21_X1 _937_ (.A(_439_),
    .B1(_053_),
    .B2(_402_),
    .ZN(_031_));
 NAND2_X1 _938_ (.A1(net57),
    .A2(net29),
    .ZN(_440_));
 OAI21_X1 _939_ (.A(_440_),
    .B1(_129_),
    .B2(net57),
    .ZN(_441_));
 NAND2_X1 _940_ (.A1(_402_),
    .A2(_441_),
    .ZN(_442_));
 OAI21_X1 _941_ (.A(_442_),
    .B1(_052_),
    .B2(_402_),
    .ZN(_032_));
 NAND2_X1 _942_ (.A1(net57),
    .A2(net30),
    .ZN(_443_));
 OAI21_X1 _943_ (.A(_443_),
    .B1(_135_),
    .B2(net57),
    .ZN(_444_));
 NAND2_X1 _944_ (.A1(_402_),
    .A2(_444_),
    .ZN(_445_));
 OAI21_X1 _945_ (.A(_445_),
    .B1(_051_),
    .B2(_402_),
    .ZN(_033_));
 NAND2_X1 _946_ (.A1(net36),
    .A2(net31),
    .ZN(_446_));
 OAI21_X1 _947_ (.A(_446_),
    .B1(_153_),
    .B2(net36),
    .ZN(_447_));
 NAND2_X1 _948_ (.A1(_402_),
    .A2(_447_),
    .ZN(_448_));
 OAI21_X1 _949_ (.A(_448_),
    .B1(_044_),
    .B2(_402_),
    .ZN(_034_));
 NAND2_X1 _950_ (.A1(net36),
    .A2(net32),
    .ZN(_449_));
 OAI21_X1 _951_ (.A(_449_),
    .B1(_170_),
    .B2(net36),
    .ZN(_450_));
 NAND2_X1 _952_ (.A1(_402_),
    .A2(_450_),
    .ZN(_451_));
 OAI21_X1 _953_ (.A(_451_),
    .B1(_043_),
    .B2(_402_),
    .ZN(_035_));
 DFF_X2 \ctrl.state.out[0]$_DFF_P_  (.D(_000_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net36),
    .QN(_003_));
 DFF_X1 \ctrl.state.out[1]$_DFF_P_  (.D(_001_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\ctrl.state.out[1] ),
    .QN(_485_));
 DFF_X1 \ctrl.state.out[2]$_DFF_P_  (.D(_002_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\ctrl.state.out[2] ),
    .QN(_484_));
 DFF_X1 \dpath.a_reg.out[0]$_DFFE_PP_  (.D(_004_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in0[0] ),
    .QN(_483_));
 DFF_X1 \dpath.a_reg.out[10]$_DFFE_PP_  (.D(_005_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in0[10] ),
    .QN(_482_));
 DFF_X1 \dpath.a_reg.out[11]$_DFFE_PP_  (.D(_006_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in0[11] ),
    .QN(_481_));
 DFF_X1 \dpath.a_reg.out[12]$_DFFE_PP_  (.D(_007_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in0[12] ),
    .QN(_480_));
 DFF_X1 \dpath.a_reg.out[13]$_DFFE_PP_  (.D(_008_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in0[13] ),
    .QN(_479_));
 DFF_X1 \dpath.a_reg.out[14]$_DFFE_PP_  (.D(_009_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in0[14] ),
    .QN(_478_));
 DFF_X1 \dpath.a_reg.out[15]$_DFFE_PP_  (.D(_010_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in0[15] ),
    .QN(_477_));
 DFF_X1 \dpath.a_reg.out[1]$_DFFE_PP_  (.D(_011_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in0[1] ),
    .QN(_476_));
 DFF_X1 \dpath.a_reg.out[2]$_DFFE_PP_  (.D(_012_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in0[2] ),
    .QN(_475_));
 DFF_X1 \dpath.a_reg.out[3]$_DFFE_PP_  (.D(_013_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in0[3] ),
    .QN(_474_));
 DFF_X1 \dpath.a_reg.out[4]$_DFFE_PP_  (.D(_014_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in0[4] ),
    .QN(_473_));
 DFF_X1 \dpath.a_reg.out[5]$_DFFE_PP_  (.D(_015_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in0[5] ),
    .QN(_472_));
 DFF_X1 \dpath.a_reg.out[6]$_DFFE_PP_  (.D(_016_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in0[6] ),
    .QN(_471_));
 DFF_X1 \dpath.a_reg.out[7]$_DFFE_PP_  (.D(_017_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in0[7] ),
    .QN(_470_));
 DFF_X1 \dpath.a_reg.out[8]$_DFFE_PP_  (.D(_018_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in0[8] ),
    .QN(_469_));
 DFF_X1 \dpath.a_reg.out[9]$_DFFE_PP_  (.D(_019_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in0[9] ),
    .QN(_468_));
 DFF_X1 \dpath.b_reg.out[0]$_DFFE_PP_  (.D(_020_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in1[0] ),
    .QN(_467_));
 DFF_X1 \dpath.b_reg.out[10]$_DFFE_PP_  (.D(_021_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in1[10] ),
    .QN(_466_));
 DFF_X1 \dpath.b_reg.out[11]$_DFFE_PP_  (.D(_022_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in1[11] ),
    .QN(_465_));
 DFF_X1 \dpath.b_reg.out[12]$_DFFE_PP_  (.D(_023_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in1[12] ),
    .QN(_464_));
 DFF_X1 \dpath.b_reg.out[13]$_DFFE_PP_  (.D(_024_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in1[13] ),
    .QN(_463_));
 DFF_X1 \dpath.b_reg.out[14]$_DFFE_PP_  (.D(_025_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in1[14] ),
    .QN(_462_));
 DFF_X1 \dpath.b_reg.out[15]$_DFFE_PP_  (.D(_026_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in1[15] ),
    .QN(_461_));
 DFF_X1 \dpath.b_reg.out[1]$_DFFE_PP_  (.D(_027_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in1[1] ),
    .QN(_460_));
 DFF_X1 \dpath.b_reg.out[2]$_DFFE_PP_  (.D(_028_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in1[2] ),
    .QN(_459_));
 DFF_X1 \dpath.b_reg.out[3]$_DFFE_PP_  (.D(_029_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in1[3] ),
    .QN(_458_));
 DFF_X1 \dpath.b_reg.out[4]$_DFFE_PP_  (.D(_030_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in1[4] ),
    .QN(_457_));
 DFF_X1 \dpath.b_reg.out[5]$_DFFE_PP_  (.D(_031_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in1[5] ),
    .QN(_456_));
 DFF_X1 \dpath.b_reg.out[6]$_DFFE_PP_  (.D(_032_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in1[6] ),
    .QN(_455_));
 DFF_X1 \dpath.b_reg.out[7]$_DFFE_PP_  (.D(_033_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in1[7] ),
    .QN(_454_));
 DFF_X1 \dpath.b_reg.out[8]$_DFFE_PP_  (.D(_034_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in1[8] ),
    .QN(_453_));
 DFF_X1 \dpath.b_reg.out[9]$_DFFE_PP_  (.D(_035_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in1[9] ),
    .QN(_452_));
 BUF_X1 input18 (.A(req_msg[25]),
    .Z(net18));
 BUF_X1 input19 (.A(req_msg[26]),
    .Z(net19));
 BUF_X1 input20 (.A(req_msg[27]),
    .Z(net20));
 BUF_X1 input21 (.A(req_msg[28]),
    .Z(net21));
 BUF_X1 input22 (.A(req_msg[29]),
    .Z(net22));
 BUF_X1 input23 (.A(req_msg[2]),
    .Z(net23));
 BUF_X1 input24 (.A(req_msg[30]),
    .Z(net24));
 BUF_X1 input25 (.A(req_msg[31]),
    .Z(net25));
 BUF_X1 input26 (.A(req_msg[3]),
    .Z(net26));
 BUF_X1 input27 (.A(req_msg[4]),
    .Z(net27));
 BUF_X1 input28 (.A(req_msg[5]),
    .Z(net28));
 BUF_X1 input29 (.A(req_msg[6]),
    .Z(net29));
 BUF_X1 input30 (.A(req_msg[7]),
    .Z(net30));
 BUF_X1 input31 (.A(req_msg[8]),
    .Z(net31));
 BUF_X1 input32 (.A(req_msg[9]),
    .Z(net32));
 BUF_X1 input33 (.A(req_val),
    .Z(net33));
 BUF_X1 input34 (.A(reset),
    .Z(net34));
 BUF_X1 input35 (.A(resp_rdy),
    .Z(net35));
 BUF_X1 output36 (.A(net57),
    .Z(req_rdy));
 BUF_X1 output37 (.A(net37),
    .Z(resp_msg[0]));
 BUF_X1 output38 (.A(net38),
    .Z(resp_msg[10]));
 BUF_X1 output39 (.A(net39),
    .Z(resp_msg[11]));
 BUF_X1 output40 (.A(net40),
    .Z(resp_msg[12]));
 BUF_X1 output41 (.A(net41),
    .Z(resp_msg[13]));
 BUF_X4 output42 (.A(net42),
    .Z(resp_msg[14]));
 BUF_X1 output43 (.A(net43),
    .Z(resp_msg[15]));
 BUF_X1 output44 (.A(net44),
    .Z(resp_msg[1]));
 BUF_X1 output45 (.A(net45),
    .Z(resp_msg[2]));
 BUF_X1 output46 (.A(net46),
    .Z(resp_msg[3]));
 BUF_X1 output47 (.A(net47),
    .Z(resp_msg[4]));
 BUF_X1 output48 (.A(net48),
    .Z(resp_msg[5]));
 BUF_X1 output49 (.A(net49),
    .Z(resp_msg[6]));
 BUF_X1 output50 (.A(net50),
    .Z(resp_msg[7]));
 BUF_X1 output51 (.A(net51),
    .Z(resp_msg[8]));
 BUF_X1 output52 (.A(net52),
    .Z(resp_msg[9]));
 BUF_X1 output53 (.A(net53),
    .Z(resp_val));
 CLKBUF_X3 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 BUF_X2 place56 (.A(_314_),
    .Z(net56));
 BUF_X4 place57 (.A(net36),
    .Z(net57));
 CLKBUF_X3 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 CLKBUF_X3 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 CLKBUF_X3 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 CLKBUF_X1 clkload0 (.A(clknet_2_0__leaf_clk));
 INV_X2 clkload1 (.A(clknet_2_1__leaf_clk));
 CLKBUF_X1 clkload2 (.A(clknet_2_2__leaf_clk));
 BUF_X1 rebuffer58 (.A(\dpath.a_lt_b$in1[11] ),
    .Z(net58));
 BUF_X1 rebuffer59 (.A(_048_),
    .Z(net59));
 BUF_X1 rebuffer60 (.A(net74),
    .Z(net60));
 BUF_X1 rebuffer61 (.A(net74),
    .Z(net61));
 BUF_X4 rebuffer62 (.A(\dpath.a_lt_b$in1[3] ),
    .Z(net62));
 BUF_X1 rebuffer63 (.A(\dpath.a_lt_b$in0[2] ),
    .Z(net63));
 BUF_X2 rebuffer64 (.A(\dpath.a_lt_b$in0[8] ),
    .Z(net64));
 BUF_X2 rebuffer65 (.A(\dpath.a_lt_b$in1[2] ),
    .Z(net65));
 BUF_X1 rebuffer66 (.A(\dpath.a_lt_b$in0[5] ),
    .Z(net66));
 BUF_X2 rebuffer67 (.A(\dpath.a_lt_b$in0[6] ),
    .Z(net67));
 BUF_X2 rebuffer68 (.A(\dpath.a_lt_b$in0[10] ),
    .Z(net68));
 BUF_X1 rebuffer69 (.A(_091_),
    .Z(net69));
 BUF_X1 rebuffer70 (.A(_248_),
    .Z(net70));
 BUF_X1 rebuffer71 (.A(_251_),
    .Z(net71));
 BUF_X1 rebuffer72 (.A(\dpath.a_lt_b$in1[8] ),
    .Z(net72));
 BUF_X1 rebuffer73 (.A(_231_),
    .Z(net73));
 BUF_X1 rebuffer74 (.A(\dpath.a_lt_b$in1[12] ),
    .Z(net74));
 BUF_X1 rebuffer75 (.A(\dpath.a_lt_b$in0[4] ),
    .Z(net75));
 BUF_X2 rebuffer76 (.A(_101_),
    .Z(net76));
 BUF_X1 rebuffer77 (.A(net114),
    .Z(net77));
 BUF_X1 rebuffer78 (.A(_098_),
    .Z(net78));
 BUF_X1 rebuffer79 (.A(_232_),
    .Z(net79));
 BUF_X1 rebuffer80 (.A(_107_),
    .Z(net80));
 BUF_X1 rebuffer81 (.A(_093_),
    .Z(net81));
 BUF_X4 rebuffer82 (.A(_121_),
    .Z(net82));
 BUF_X1 rebuffer83 (.A(_274_),
    .Z(net83));
 BUF_X1 rebuffer84 (.A(_159_),
    .Z(net84));
 BUF_X1 rebuffer85 (.A(_074_),
    .Z(net85));
 BUF_X1 rebuffer86 (.A(net125),
    .Z(net86));
 BUF_X4 rebuffer87 (.A(_134_),
    .Z(net87));
 BUF_X4 rebuffer88 (.A(_107_),
    .Z(net88));
 BUF_X1 rebuffer89 (.A(\dpath.a_lt_b$in1[13] ),
    .Z(net89));
 BUF_X1 rebuffer91 (.A(_255_),
    .Z(net91));
 BUF_X1 rebuffer110 (.A(net51),
    .Z(net110));
 BUF_X4 rebuffer111 (.A(_151_),
    .Z(net111));
 BUF_X1 rebuffer113 (.A(\dpath.a_lt_b$in1[6] ),
    .Z(net113));
 BUF_X1 rebuffer114 (.A(_089_),
    .Z(net114));
 BUF_X1 rebuffer115 (.A(\dpath.a_lt_b$in1[7] ),
    .Z(net115));
 BUF_X1 rebuffer125 (.A(_227_),
    .Z(net125));
 BUF_X1 rebuffer126 (.A(_249_),
    .Z(net126));
 BUF_X2 rebuffer127 (.A(\dpath.a_lt_b$in0[14] ),
    .Z(net127));
 BUF_X1 rebuffer128 (.A(_273_),
    .Z(net128));
 BUF_X4 rebuffer132 (.A(\dpath.a_lt_b$in0[4] ),
    .Z(net132));
 BUF_X1 rebuffer133 (.A(net50),
    .Z(net133));
 BUF_X2 rebuffer134 (.A(_151_),
    .Z(net134));
 BUF_X1 rebuffer137 (.A(net38),
    .Z(net137));
 NAND2_X4 clone138 (.A1(_297_),
    .A2(_304_),
    .ZN(net138));
 BUF_X2 rebuffer139 (.A(_081_),
    .Z(net139));
 NAND4_X2 clone141 (.A1(_297_),
    .A2(\ctrl.state.out[2] ),
    .A3(_003_),
    .A4(_304_),
    .ZN(net141));
 BUF_X2 rebuffer143 (.A(\dpath.a_lt_b$in0[7] ),
    .Z(net143));
endmodule
